CPU_FSM.bsv