package DUT;

String title   = "The C Programming Language";
String authors = "Kernighan and Ritchie";

Bit #(11) year = 1978;

Bit #(4)  month = 2;

Bit #(5)  day = 22;

endpackage
