module mkTop (Empty);

   rule rl_once;
      $display ("Hello, World!");
      $finish (0);
   endrule

endmodule
